`timescale 1ns / 1ps

module ForwardingControl(Instruction_EX,RegDst_MEM,Reg_Dst_WB,ALUResult_MEM,RegData_WB,ReadData1Sel,ReadData2Sel);
	input [31:0] Instruction_EX,ALUResult_MEM;
	
	
	
endmodule